//Este modulo controla los datos enviados a los puertos del display

module module_display #(

    input logic [3 : 0] binary_code,     //Entrada: Código Grey ya convertido a binario
    output logic [6 : 0] display_code
);

endmodule