//Este módulo interconecta los tres sub módulos 