//Este modulo codifica BCD a 7 segmentos 