//Este modulo controla los datos enviados a los puertos del display

module display #(

    input logic [3 : 0] binary_code,     
    output logic [6 : 0] display_code



);

endmodule